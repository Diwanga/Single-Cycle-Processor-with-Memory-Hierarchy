//////////////////////////////////////////////////////////////////
//module for making two's compliment
//////////////////////////////////////////////////////////////////

module compliment(OUT,IN);   
output [7:0] OUT;
input [7:0] IN;

assign OUT= ~IN+1'b1;  //making two's compliment of input 

endmodule





///////////////////////////////////////////////////////////////////////////////////////

